library IEEE;
use IEEE.std_logic_1164.all;

entity decoder_5_32 is

  port(sel       : in std_logic_vector(4 downto 0);
       wr	 : in std_logic;
       output    : out std_logic_vector(31 downto 0));

end decoder_5_32;

architecture dataflow of decoder_5_32 is


begin

output <= "00000000000000000000000000000001" when sel = "00000" and wr='1' else 
"00000000000000000000000000000010" when sel = "00001" and wr='1' else 
"00000000000000000000000000000100" when sel = "00010" and wr='1' else 
"00000000000000000000000000001000" when sel = "00011" and wr='1' else 
"00000000000000000000000000010000" when sel = "00100" and wr='1' else 
"00000000000000000000000000100000" when sel = "00101" and wr='1' else 
"00000000000000000000000001000000" when sel = "00110" and wr='1' else 
"00000000000000000000000010000000" when sel = "00111" and wr='1' else 
"00000000000000000000000100000000" when sel = "01000" and wr='1' else
"00000000000000000000001000000000" when sel = "01001" and wr='1' else
"00000000000000000000010000000000" when sel = "01010" and wr='1' else
"00000000000000000000100000000000" when sel = "01011" and wr='1' else
"00000000000000000001000000000000" when sel = "01100" and wr='1' else
"00000000000000000010000000000000" when sel = "01101" and wr='1' else
"00000000000000000100000000000000" when sel = "01110" and wr='1' else
"00000000000000001000000000000000" when sel = "01111" and wr='1' else
"00000000000000010000000000000000" when sel = "10000" and wr='1' else
"00000000000000100000000000000000" when sel = "10001" and wr='1' else
"00000000000001000000000000000000" when sel = "10010" and wr='1' else
"00000000000010000000000000000000" when sel = "10011" and wr='1' else
"00000000000100000000000000000000" when sel = "10100" and wr='1' else
"00000000001000000000000000000000" when sel = "10101" and wr='1' else
"00000000010000000000000000000000" when sel = "10110" and wr='1' else
"00000000100000000000000000000000" when sel = "10111" and wr='1' else
"00000001000000000000000000000000" when sel = "11000" and wr='1' else
"00000010000000000000000000000000" when sel = "11001" and wr='1' else
"00000100000000000000000000000000" when sel = "11010" and wr='1' else
"00001000000000000000000000000000" when sel = "11011" and wr='1' else
"00010000000000000000000000000000" when sel = "11100" and wr='1' else
"00100000000000000000000000000000" when sel = "11101" and wr='1' else
"01000000000000000000000000000000" when sel = "11110" and wr='1' else
"10000000000000000000000000000000" when sel = "11111" and wr='1' else
"00000000000000000000000000000000";

end dataflow;